module and_gate_tb;
    reg a, b;
    wire y;
    and_gate dut (
           .a1(a),
           .b1(b),
           .y1(y)
    );
   initial begin
      $dumpfile("and_gate.vcd");
      $dumpvars(0, and_gate_tb);
      $monitor("Time=%0t | a=%b b=%b | y=%b", $time, a, b, y);
      a = 0; b = 0;
      #10 a = 0; b = 1;
      #10 a = 1; b = 0;
      #10 a = 1; b = 1;
      #10;
      $finish;
   end
endmodule
  

