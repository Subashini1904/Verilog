module d_ff_sync_rst (
input clk,
input rst,      
input d,
output reg q
);
always @(posedge clk) begin
    if (rst)
        q <= 1'b0;   
    else
        q <= d;
end
endmodule


//OUTPUT//
Time  clk  rst  d  q
0    0     1    0  x
3    0     0    0  x
5    1     0    0  0
7    1     0    1  0
10    0    0    1  0
13    0    0    0  0
15    1    1    0  0
19    1    0    0  0
20    0    0    0  0
25    1    0    0  0
30    0    0    0  0
35    1    0    0  0
