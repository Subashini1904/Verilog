module andgate_if_tb;
reg a,b;
wire y;
andgate_if dut(
.a(a),
.b(b),
.y(y)
);
initial begin
  $dumpfile("andgate_if.vcd");
  $dumpvars(0, andgate_if_tb);
  $monitor("time=%0t | a=%b b=%b | y=%b", $time, a, b, y);
  a=0;b=0;#10;
  a=0;b=1;#10;
  a=1;b=0;#10;
  a=1;b=1;#10;
  $finish;
  end
endmodule
