module mux16to1_4to1 (
input  [15:0] in,
input  [3:0]  s,
output y
);
wire w0, w1, w2, w3;
assign w0 = (s[1:0] == 2'b00) ? in[0]:
            (s[1:0] == 2'b01) ? in[1]:
            (s[1:0] == 2'b10) ? in[2]:
                                in[3];
assign w1 = (s[1:0] == 2'b00) ? in[4]:
            (s[1:0] == 2'b01) ? in[5]:
            (s[1:0] == 2'b10) ? in[6]:
                                in[7];
assign w2 = (s[1:0] == 2'b00) ? in[8]:
            (s[1:0] == 2'b01) ? in[9]:
            (s[1:0] == 2'b10) ? in[10]:
                                in[11];
assign w3 = (s[1:0] == 2'b00) ? in[12]:
            (s[1:0] == 2'b01) ? in[13]:
            (s[1:0] == 2'b10) ? in[14]:
                                in[15];
assign y = (s[3:2] == 2'b00) ? w0:
           (s[3:2] == 2'b01) ? w1:
           (s[3:2] == 2'b10) ? w2:
                               w3;

endmodule


//OUTPUT//
time=0 | in=1010110001101001 | s=0 | y=1
time=10 | in=1010110001101001 | s=1 | y=0
time=20 | in=1010110001101001 | s=2 | y=0
time=30 | in=1010110001101001 | s=3 | y=1
time=40 | in=1010110001101001 | s=4 | y=0
time=50 | in=1010110001101001 | s=5 | y=1
time=60 | in=1010110001101001 | s=6 | y=1
time=70 | in=1010110001101001 | s=7 | y=0
time=80 | in=1010110001101001 | s=8 | y=0
time=90 | in=1010110001101001 | s=9 | y=0
time=100 | in=1010110001101001 | s=10 | y=1
time=110 | in=1010110001101001 | s=11 | y=1
time=120 | in=1010110001101001 | s=12 | y=0
time=130 | in=1010110001101001 | s=13 | y=1
time=140 | in=1010110001101001 | s=14 | y=0
time=150 | in=1010110001101001 | s=15 | y=1
