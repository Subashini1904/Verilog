module and_gate(input a1, b1, output y1);
   assign y1 = a1 & b1;
endmodule
 
